`define MAC_SOURCE_REPLACE_EN 1
`define MAC_TARGET_CHECK_EN 1
`define MAC_BROADCAST_FILTER_EN 1
`define MAC_TX_FF_DEPTH 9
`define MAC_RX_FF_DEPTH 9
`define MAC_TARGET_XILINX 1
// `define MAC_TARGET_ALTERA 1
