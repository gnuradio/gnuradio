
module traffic_cop();


endmodule // traffic_cop



/*
 
 Traffic Cop to control buffer pool
 
 Inputs
 
 Commands
 
 Basic Operations
 
 Outputs
 
 
 
 
 
 */
