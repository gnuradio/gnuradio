module xlnx_glbl
(
  GSR,
  GTS
);

  //--------------------------------------------------------------------------
  // Parameters
  //--------------------------------------------------------------------------

  //--------------------------------------------------------------------------
  // IO declarations
  //--------------------------------------------------------------------------

  output GSR;
  output GTS;

  //--------------------------------------------------------------------------
  // Local declarations
  //--------------------------------------------------------------------------

  //--------------------------------------------------------------------------
  // Internal declarations
  //--------------------------------------------------------------------------

  assign GSR = 0;
  assign GTS = 0;
  
endmodule
