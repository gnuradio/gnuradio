-------------------------------------------------------------------------------
--
-- SD/MMC Bootloader
--
-- $Id: spi_counter-c.vhd,v 1.1 2005/02/08 20:41:33 arniml Exp $
--
-------------------------------------------------------------------------------

configuration spi_counter_rtl_c0 of spi_counter is

  for rtl
  end for;

end spi_counter_rtl_c0;
